package types_pkg;

typedef struct packed {logic a, b, c;} input_signals_t;
typedef struct packed {logic x, y, z;} output_signals_t;
typedef struct packed {logic [2:0] params;} parameters_t;

endpackage
