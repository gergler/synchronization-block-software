module freDetect(clk, test, rst, q);  
  input clk;
  input test; 
  input rst; 
	
  wire count_en;
  wire latch_en;
  wire clear;

  output[31:0] q;

  control u_control(.clk(clk), .rst(rst), .count_en(count_en), .latch_en(latch_en), .clear(clear));  
  counter u_counter(.count_en(count_en), .clear(clear), .rst(rst), .test(test), .q(q)); 
     
endmodule  

module control(clk, rst, count_en, latch_en, clear);  

  input clk;  
  input rst;  
  output count_en;  
  output latch_en;  
  output clear;  

  reg[1:0] state; // \u0421\u0438\u0433\u043d\u0430\u043b \u0441\u043e\u0441\u0442\u043e\u044f\u043d\u0438\u044f, \u0438\u0441\u043f\u043e\u043b\u044c\u0437\u0443\u0435\u043c\u044b\u0439 \u0434\u043b\u044f \u0443\u043f\u0440\u0430\u0432\u043b\u0435\u043d\u0438\u044f \u0440\u0430\u0437\u043b\u0438\u0447\u043d\u044b\u043c\u0438 \u0441\u0438\u0433\u043d\u0430\u043b\u0430\u043c\u0438 \u0432\u043a\u043b\u044e\u0447\u0435\u043d\u0438\u044f  
  reg count_en;  
  reg latch_en;  
  reg clear;  

  always @(posedge clk or negedge rst)  
  if(!rst) // \u0421\u0438\u0433\u043d\u0430\u043b \u0441\u0431\u0440\u043e\u0441\u0430 \u0434\u0435\u0439\u0441\u0442\u0432\u0438\u0442\u0435\u043b\u0435\u043d  
    begin  // \u0423\u0434\u0430\u043b\u044f\u0435\u043c \u0440\u0430\u0437\u043b\u0438\u0447\u043d\u044b\u0435 \u0440\u0430\u0437\u0440\u0435\u0448\u0430\u044e\u0449\u0438\u0435 \u0441\u0438\u0433\u043d\u0430\u043b\u044b  
      state <= 2'd0;  
      count_en <= 1'b0;  
      latch_en <=1'b0;  
      clear <= 1'b0;  
    end  
   else 
      	2'd0:   
          begin // \u041f\u0435\u0440\u0432\u044b\u0439 \u043f\u0435\u0440\u0435\u0434\u043d\u0438\u0439 \u0444\u0440\u043e\u043d\u0442 \u043f\u0440\u0438\u0445\u043e\u0434\u0438\u0442, \u043d\u0430\u0447\u0430\u0442\u044c \u043f\u043e\u0434\u0441\u0447\u0435\u0442, \u043f\u043e\u0434\u0441\u0447\u0438\u0442\u0430\u0442\u044c \u0447\u0438\u0441\u043b\u043e \u043d\u0430\u0440\u0430\u0441\u0442\u0430\u044e\u0449\u0438\u0445 \u0444\u0440\u043e\u043d\u0442\u043e\u0432 \u0441\u0438\u0433\u043d\u0430\u043b\u0430 \u043f\u0440\u0438 \u0438\u0441\u043f\u044b\u0442\u0430\u043d\u0438\u0438 \u0432 \u0442\u0435\u0447\u0435\u043d\u0438\u0435 1 \u043e\u043f\u043e\u0440\u043d\u043e\u0433\u043e \u0441\u0438\u0433\u043d\u0430\u043b\u0430, \u044d\u0442\u043e \u0447\u0438\u0441\u043b\u043e \u044f\u0432\u043b\u044f\u0435\u0442\u0441\u044f \u0447\u0430\u0441\u0442\u043e\u0442\u0430 \u0441\u0438\u0433\u043d\u0430\u043b\u0430 \u043f\u0440\u0438 \u0438\u0441\u043f\u044b\u0442\u0430\u043d\u0438\u0438  
            count_en <= 1'b1;  // \u0421\u0438\u0433\u043d\u0430\u043b \u0432\u043a\u043b\u044e\u0447\u0435\u043d\u0438\u044f \u043f\u043e\u0434\u0441\u0447\u0435\u0442\u0430 \u0434\u0435\u0439\u0441\u0442\u0432\u0438\u0442\u0435\u043b\u0435\u043d  
            latch_en <=1'b0;  
            clear <= 1'b0;  
            state <= 2'd1;  
          end  
        2'd1:  
          begin // \u041f\u0440\u0438\u0445\u043e\u0434\u0438\u0442 \u0432\u0442\u043e\u0440\u043e\u0439 \u043d\u0430\u0440\u0430\u0441\u0442\u0430\u044e\u0449\u0438\u0439 \u0444\u0440\u043e\u043d\u0442, \u0441\u0447\u0435\u0442 \u0437\u0430\u0432\u0435\u0440\u0448\u0435\u043d, \u0441\u0438\u0433\u043d\u0430\u043b \u0440\u0430\u0437\u0440\u0435\u0448\u0435\u043d\u0438\u044f \u0444\u0438\u043a\u0441\u0430\u0446\u0438\u0438 \u0434\u0435\u0439\u0441\u0442\u0432\u0438\u0442\u0435\u043b\u0435\u043d, \u0438 \u0438\u0437\u043c\u0435\u0440\u0435\u043d\u043d\u0430\u044f \u0447\u0430\u0441\u0442\u043e\u0442\u0430 \u0444\u0438\u043a\u0441\u0438\u0440\u0443\u0435\u0442\u0441\u044f \u0432 \u0437\u0430\u0449\u0435\u043b\u043a\u0435  
            count_en <= 1'b0;  
            latch_en <=1'b1;  
            clear <= 1'b0;  
            state <= 2'd2;  
          end  
        2'd2:   
          begin // \u041f\u043e\u044f\u0432\u043b\u044f\u0435\u0442\u0441\u044f \u0442\u0440\u0435\u0442\u0438\u0439 \u043d\u0430\u0440\u0430\u0441\u0442\u0430\u044e\u0449\u0438\u0439 \u0444\u0440\u043e\u043d\u0442, \u0441\u0438\u0433\u043d\u0430\u043b \u0440\u0430\u0437\u0440\u0435\u0448\u0435\u043d\u0438\u044f \u0441\u0431\u0440\u043e\u0441\u0430 \u0434\u0435\u0439\u0441\u0442\u0432\u0438\u0442\u0435\u043b\u0435\u043d, \u0438 \u0441\u0447\u0435\u0442\u0447\u0438\u043a \u043e\u0447\u0438\u0449\u0430\u0435\u0442\u0441\u044f \u0434\u043b\u044f \u043f\u043e\u0434\u0433\u043e\u0442\u043e\u0432\u043a\u0438 \u043a \u0441\u043b\u0435\u0434\u0443\u044e\u0449\u0435\u043c\u0443 \u0441\u0447\u0435\u0442\u0443  
            count_en <= 1'b0;  
            latch_en <=1'b0;  
            clear <= 1'b1;  
            state <= 2'd0; // \u0421\u043e\u0441\u0442\u043e\u044f\u043d\u0438\u0435 \u043e\u0447\u0438\u0449\u0430\u0435\u0442\u0441\u044f \u0438 \u043f\u0435\u0440\u0435\u0445\u043e\u0434\u0438\u043c \u043a \u0441\u043b\u0435\u0434\u0443\u044e\u0449\u0435\u043c\u0443 \u0438\u0437\u043c\u0435\u0440\u0435\u043d\u0438\u044e  
          end  
        default:  
          begin  
            count_en <= 1'b0;  
            latch_en <=1'b0;  
            clear <= 1'b0;  
            state <= 2'd0;  
          end          
      endcase             
    end      
endmodule  
  
// \u041c\u043e\u0434\u0443\u043b\u044c \u043f\u043e\u0434\u0441\u0447\u0435\u0442\u0430  
module counter(count_en, rst, clear, test, q);  
  input count_en;
  input rst;   // \u0421\u0431\u0440\u043e\u0441 \u0441\u0438\u0433\u043d\u0430\u043b\u0430  
  input clear; // \u041e\u0447\u0438\u0441\u0442\u0438\u0442\u044c \u0441\u0438\u0433\u043d\u0430\u043b  
  input test;   // \u0421\u0438\u0433\u043d\u0430\u043b \u0434\u043b\u044f \u0442\u0435\u0441\u0442\u0438\u0440\u043e\u0432\u0430\u043d\u0438\u044f    
  output reg[31:0] q;
    
  always @(posedge test or negedge rst) // \u0412\u0432\u043e\u0434 \u043d\u0430\u0440\u0430\u0441\u0442\u0430\u044e\u0449\u0435\u0433\u043e \u0444\u0440\u043e\u043d\u0442\u0430 \u0438\u0437\u043c\u0435\u0440\u044f\u0435\u043c\u043e\u0433\u043e \u0441\u0438\u0433\u043d\u0430\u043b\u0430 \u043a\u0430\u043a \u0447\u0443\u0432\u0441\u0442\u0432\u0438\u0442\u0435\u043b\u044c\u043d\u043e\u0433\u043e \u0441\u0438\u0433\u043d\u0430\u043b\u0430  
  if(!rst) // \u0421\u0438\u0433\u043d\u0430\u043b \u0441\u0431\u0440\u043e\u0441\u0430 \u0434\u0435\u0439\u0441\u0442\u0432\u0438\u0442\u0435\u043b\u0435\u043d, \u0438 \u0432\u044b\u0445\u043e\u0434 \u0441\u0447\u0435\u0442\u0447\u0438\u043a\u0430 \u043e\u0447\u0438\u0449\u0430\u0435\u0442\u0441\u044f  
      begin  
        q <= 0;  
      end  
        
  else if(count_en) // \u0421\u0438\u0433\u043d\u0430\u043b \u0440\u0430\u0437\u0440\u0435\u0448\u0435\u043d\u0438\u044f \u043f\u043e\u0434\u0441\u0447\u0435\u0442\u0430
      begin // q \u0443\u0432\u0435\u043b\u0438\u0447\u0438\u0432\u0430\u0435\u0442\u0441\u044f \u043d\u0430 1 \u043a\u0430\u0436\u0434\u044b\u0439 \u0440\u0430\u0437, \u043a\u043e\u0433\u0434\u0430 \u0434\u043e\u0441\u0442\u0438\u0433\u0430\u0435\u0442\u0441\u044f \u043d\u0430\u0440\u0430\u0441\u0442\u0430\u044e\u0449\u0438\u0439 \u0444\u0440\u043e\u043d\u0442 \u0438\u0437\u043c\u0435\u0440\u044f\u0435\u043c\u043e\u0433\u043e \u0441\u0438\u0433\u043d\u0430\u043b\u0430  
          begin  
            q <= q + 1;
	    $display("period/clk = %b", q);
          end  
      end  
        
   else if(clear) // \u0415\u0441\u043b\u0438 \u0441\u0438\u0433\u043d\u0430\u043b \u043e\u0447\u0438\u0441\u0442\u043a\u0438 \u0434\u0435\u0439\u0441\u0442\u0432\u0438\u0442\u0435\u043b\u0435\u043d, \u0441\u0447\u0435\u0442\u0447\u0438\u043a \u043e\u0447\u0438\u0449\u0430\u0435\u0442\u0441\u044f, \u0432 \u043e\u0441\u043d\u043e\u0432\u043d\u043e\u043c \u0438\u0441\u043f\u043e\u043b\u044c\u0437\u0443\u0435\u0442\u0441\u044f \u0434\u043b\u044f \u043f\u043e\u0434\u0433\u043e\u0442\u043e\u0432\u043a\u0438 \u043a \u0441\u043b\u0435\u0434\u0443\u044e\u0449\u0435\u043c\u0443 \u0438\u0437\u043c\u0435\u0440\u0435\u043d\u0438\u044e  
      	begin  
          q <= 0;  
      	end  

   else  
   	begin  
    	  q <= q;  
    	end   
    
endmodule  